module  ID_EX_PipelineReg (
    input clk, rst_n, ReadIn, WriteReg, PCS, MemtoReg, MemRead, MemWrite, B, BR, HLT,
    input [1:0] AluSrc1, AluSrc2,
    input [2:0] AluOp,
    input [15:0] ReadData1, ReadData2
);

//Excute Stage Signals


//Memory Stage Signals

//Write Back Stage Signals

//
    
endmodule